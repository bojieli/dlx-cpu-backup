module main();
endmodule // main
